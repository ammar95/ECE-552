module cache_tb();

